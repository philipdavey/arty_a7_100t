------------------------------------------------------------------------------
-- Title       :
-- Project     : 
------------------------------------------------------------------------------
-- File        :
-- Author      :
------------------------------------------------------------------------------
-- Description :
------------------------------------------------------------------------------

------------------------------------------------------------------------------
-- Library declaration :
------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

------------------------------------------------------------------------------
-- Entity declaration :
------------------------------------------------------------------------------
entity arty_top is
  port (
    fpga_clk_100_mhz : std_logic;
    fpga_rst_n       : std_logic
  );
end arty_top;

------------------------------------------------------------------------------
-- Architecture declaration :
------------------------------------------------------------------------------
architecture rtl_arty_top of arty_top is

begin

end rtl_arty_top;